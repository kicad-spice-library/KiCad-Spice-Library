Test file for the 'alter' command

.model BC107    NPN(Is=1.527f Xti=3 Eg=1.11 Vaf=106.8 Bf=334.5 Ne=1.642
+               Ise=222f Ikf=.1596 Xtb=1.5 Br=.788 Nc=2 Isc=0 Ikr=0 Re=.6 Rc=0.25
+               Cjc=6.072p Mjc=.3333 Vjc=.75 Fc=.5 Cje=10.67p Mje=.3333 Vje=.75
+               Tr=10n Tf=471.8p Itf=0 Vtf=0 Xtf=0)

* Circuit to plot curves of Ic versus Vce for comparison with a datasheet

Ib 0 base DC 50e-6

*  C B E model
Q1 collector base emitter BC107

Rc collector 10 10k
Re emitter   0  1k

Vce 10 0 10V

*#op
*#print base collector emitter vce#branch v(10)

* -- BJT instance output
*#print @q1[off] @q1[icvbe] @q1[icvce] @q1[area] @q1[temp]
*#print @q1[colnode] @q1[basenode] @q1[emitnode] @q1[substnode] @q1[colprimenode] @q1[emitprimenode]
*#print @q1[ic]
*#print @q1[ib]
*#print @q1[ie]
*#print @q1[is]
*#print @q1[vbe] @q1[vbc] @q1[gm] @q1[gpi] @q1[gmu] @q1[gx] @q1[go] @q1[geqcb] @q1[gccs] @q1[geqbx]
*#print @q1[cpi] @q1[cmu] @q1[cbx] @q1[ccs] @q1[cqbe] @q1[cqbc] @q1[cqcs] @q1[cqbx] @q1[cexbc]
*#print @q1[qbe] @q1[qbc] @q1[qcs] @q1[qbx] @q1[p]

* -- BJT model output
*#print @bc107[npn] @BC107[pnp] @BC107[is] @BC107[bf] @BC107[nf] @BC107[vaf] @BC107[va] @BC107[ikf]
*#print @BC107[ik] @BC107[ise] @BC107[ne] @BC107[br] @BC107[nr] @BC107[var] @BC107[vb] @BC107[ikr]
*#print @BC107[isc] @BC107[nc] @BC107[rb] @BC107[irb] @BC107[rbm] @BC107[re] @BC107[rc] @BC107[cje]
*#print @BC107[vje] @BC107[pe] @BC107[mje] @BC107[me] @BC107[tf] @BC107[xtf] @BC107[vtf] @BC107[itf]
*#print @BC107[ptf] @BC107[cjc] @BC107[vjc] @BC107[pc] @BC107[mjc] @BC107[mc] @BC107[xcjc] @BC107[tr]
*#print @BC107[cjs] @BC107[ccs] @BC107[vjs] @BC107[ps] @BC107[mjs] @BC107[ms] @BC107[xtb] @BC107[eg]
*#print @BC107[xti] @BC107[fc] @BC107[tnom] @BC107[kf] @BC107[af]
*#print @BC107[type]
*#print @BC107[invearlyvoltf] @BC107[invearlyvoltr] @BC107[invrolloffr] @BC107[collectorconduct]
*#print @BC107[emitterconduct] @BC107[transtimevbcfact] @BC107[excessphasefactor]

* -- BJT instance input
*#alter @q1[ic] = [ 0 0 ]
*#alter @q1[off] = 0
*#alter @q1[icvbe] = 0
*#alter @q1[icvce] = 0
*#alter @q1[area] = 0
*#alter @q1[temp] = 0

* -- BJT model input
*#alter @bc107[npn] = 0
*#alter @BC107[pnp] = 0
*#alter @BC107[is] = 0
*#alter @BC107[bf] = 0
*#alter @BC107[nf] = 0
*#alter @BC107[vaf] = 0
*#alter @BC107[va] = 0
*#alter @BC107[ikf] = 0
*#alter @BC107[ik] = 0
*#alter @BC107[ise] = 0
*#alter @BC107[ne] = 0
*#alter @BC107[br] = 0
*#alter @BC107[nr] = 0
*#alter @BC107[var] = 0
*#alter @BC107[vb] = 0
*#alter @BC107[ikr] = 0
*#alter @BC107[isc] = 0
*#alter @BC107[nc] = 0
*#alter @BC107[rb] = 0
*#alter @BC107[irb] = 0
*#alter @BC107[rbm] = 0
*#alter @BC107[re] = 0
*#alter @BC107[rc] = 0
*#alter @BC107[cje] = 0
*#alter @BC107[vje] = 0
*#alter @BC107[pe] = 0
*#alter @BC107[mje] = 0
*#alter @BC107[me] = 0
*#alter @BC107[tf] = 0
*#alter @BC107[xtf] = 0
*#alter @BC107[vtf] = 0
*#alter @BC107[itf] = 0
*#alter @BC107[ptf] = 0
*#alter @BC107[cjc] = 0
*#alter @BC107[vjc] = 0
*#alter @BC107[pc] = 0
*#alter @BC107[mjc] = 0
*#alter @BC107[mc] = 0
*#alter @BC107[xcjc] = 0
*#alter @BC107[tr] = 0
*#alter @BC107[cjs] = 0
*#alter @BC107[ccs] = 0
*#alter @BC107[vjs] = 0
*#alter @BC107[ps] = 0
*#alter @BC107[mjs] = 0
*#alter @BC107[ms] = 0
*#alter @BC107[xtb] = 0
*#alter @BC107[eg] = 0
*#alter @BC107[xti] = 0
*#alter @BC107[fc] = 0
*#alter @BC107[tnom] = 0
*#alter @BC107[kf] = 0
*#alter @BC107[af] = 0

* -- This should fail
*#alter @BC107[invearlyvoltf] = 0

