* Version 2.0 Copyright � Linear Technology Corp. 10/19/05. All rights reserved.
* NODES 1 AND 8 = COMPENSATION PINS
*
.SUBCKT LM101A 3 2 7 4 6 1 8 ; IN+ IN- VCC VEE OUT COMP1 COMP2
* USE C=30 PF IN MAIN CIRCUIT (CA TO CB).
* INPUT
RC1 7 80 5.895E+03
RC2 7 90 5.895E+03
Q1 80 2 10 QM1
Q2 90 3 11 QM2
C1 80 90 5.460E-12
RE1 10 12 2.438E+03
RE2 11 12 2.438E+03
IEE 12 4 1.506E-05
RE 12 0 1.328E+07
CE 12 0 1.579E-12
* INTERMEDIATE
GCM 0 8 12 0 2.689E-09
GA 8 0 80 90 1.696E-04
R2 8 0 1.000E+05
* EXTERNAL COMP CAP USED FOR C2 (SEE NOTE ABOVE).
GB 1 0 8 0 1.401E+02
* OUTPUT
RO1 1 6 3.333E+01
RO2 1 0 6.667E+01
RC 17 0 4.758E-05
GC 0 17 6 0 2.102E+04
D1 1 17 DM1
D2 17 1 DM1
D3 6 13 DM2
D4 14 6 DM2
VC 7 13 1.808E+00
VE 14 4 1.808E+00
IP 7 4 1.785E-03
DSUB 4 7 DM2
* MODELS
.MODEL QM1 NPN (IS=8.000E-16 BF=2.439E+02)
.MODEL QM2 NPN (IS=8.220E-16 BF=2.564E+02)
.MODEL DM1 D (IS=3.337E-15)
.MODEL DM2 D (IS=8.000E-16)
.ENDS LM101A
