.MODEL 20ets12a+3s d
+IS=2.797e-10 RS=0.0113232 N=1.38813 EG=1.07556
+XTI=4 BV=1200 IBV=0.0001 CJO=1e-11
+VJ=0.7 M=0.5 FC=0.5 TT=1e-09
+KF=0 AF=1
* Model generated on Apr 26, 96
* Model format: SPICE3

