Basic RC circuit
r 1 2 1.0
*l 1 2 1.0
c 2 0 1.0
vin 1 0  pulse (0 1) ac 1
.tran  0.1 7.0
*.ac dec 10 .01 10
.plot tran  v(2) i(vin)
*.plot ac  vdb(2) xlog
.end
