*MC33071 OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
*CONNECTIONS: 1=+In, 2=-In, 3=+V, 4=-V, 5=Out
.SUBCKT MC33071  1 2 3 4 5
  C1   11 12 8.660E-12
  C2    6  7 8.000E-12
  CEE  10 99 1.231E-12
  DC    5 53 DX
  DE   54  5 DX
  DLP  90 91 DX
  DLN  92 90 DX
  DP    4  3 DX
  EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
  FB    7 99 POLY(5) VB VC VE VLP VLN 0 8.842E6 
  + -9E6 9E6 9E6 -9E6
  GA    6  0 11 12 251.3E-6
  GCM   0  6 10 99 3.550E-9
  IEE   3 10 DC 120.2E-6
  HLIM 90  0 VLIM 1K
  Q1   11  2 13 QX
  Q2   12  1 14 QX
  R2    6  9 100.0E3
  RC1   4 11 3.979E3
  RC2   4 12 3.979E3
  RE1  13 10 3.542E3
  RE2  14 10 3.542E3
  REE  10 99 1.664E6
  RO1   8  5 30
  RO2   7 99 45
  RP    3  4 34.09E3
  VB    9  0 DC 0
  VC    3 53 DC 1
  VE   54  4 DC .3
  VLIM  7  8 DC 0
  VLP  91  0 DC 30
  VLN   0 92 DC 30
.MODEL DX D(IS=800.0E-18)
.MODEL QX PNP(IS=800.0E-18 BF=600)
.ENDS MC33071
 
