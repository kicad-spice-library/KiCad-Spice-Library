.MODEL 15clq100 d
+IS=6.44968e-05 RS=0.014091 N=2 EG=0.996757
+XTI=0.5 BV=100 IBV=0.005 CJO=1.38463e-09
+VJ=0.4 M=0.466344 FC=0.5 TT=0
+KF=0 AF=1
* Model generated on May 28, 96
* Model format: SPICE3

