* LM324LV - Rev. A
* Created by Paul Goedeke; June 06, 2018
* Created with Green-Williams-Lis Op Amp Macro-model Architecture
* Copyright 2018 by Texas Instruments Corporation
******************************************************
* MACRO-MODEL SIMULATED PARAMETERS:
******************************************************
* OPEN-LOOP GAIN AND PHASE VS. FREQUENCY  WITH RL, CL EFFECTS (Aol)
* UNITY GAIN BANDWIDTH (GBW)
* INPUT COMMON-MODE REJECTION RATIO VS. FREQUENCY (CMRR)
* POWER SUPPLY REJECTION RATIO VS. FREQUENCY (PSRR)
* DIFFERENTIAL INPUT IMPEDANCE (Zid)
* COMMON-MODE INPUT IMPEDANCE (Zic)
* OPEN-LOOP OUTPUT IMPEDANCE VS. FREQUENCY (Zo)
* OUTPUT CURRENT THROUGH THE SUPPLY (Iout)
* INPUT VOLTAGE NOISE DENSITY VS. FREQUENCY (en)
* INPUT CURRENT NOISE DENSITY VS. FREQUENCY (in)
* OUTPUT VOLTAGE SWING vs. OUTPUT CURRENT (Vo)
* SHORT-CIRCUIT OUTPUT CURRENT (Isc)
* QUIESCENT CURRENT (Iq)
* SETTLING TIME VS. CAPACITIVE LOAD (ts)
* SLEW RATE (SR)
* SMALL SIGNAL OVERSHOOT VS. CAPACITIVE LOAD
* LARGE SIGNAL RESPONSE
* OVERLOAD RECOVERY TIME (tor)
* INPUT BIAS CURRENT (Ib)
* INPUT OFFSET CURRENT (Ios)
* INPUT OFFSET VOLTAGE (Vos)
* INPUT COMMON-MODE VOLTAGE RANGE (Vcm)
* INPUT/OUTPUT ESD CELLS (ESDin, ESDout)
******************************************************
.subckt LM324LV IN+ IN- VCC VEE OUT
******************************************************
* MODEL DEFINITIONS:
.model BB_SW VSWITCH(Ron=50 Roff=1e12 Von=700e-3 Voff=0)
.model ESD_SW VSWITCH(Ron=50 Roff=1e12 Von=250e-3 Voff=0)
.model OL_SW VSWITCH(Ron=1e-3 Roff=1e9 Von=900e-3 Voff=800e-3)
.model OR_SW VSWITCH(Ron=10e-3 Roff=1e9 Von=1e-3 Voff=0)
*.model R_NOISELESS RES(T_ABS=-273.15)
******************************************************

I_OS        ESDn MID 7P
I_B         31 MID 10P
V_GRp       56 MID 195
V_GRn       57 MID -195
V_ISCp      50 MID 40
V_ISCn      51 MID -40
V_ORn       39 VCLP -1.45
V11         55 38 0
V_ORp       37 VCLP 1.5
V12         54 36 0
V4          27 OUT 0
VCM_MIN     77 VEE_B -100M
VCM_MAX     78 VCC_B -1.5
I_Q         VCC VEE 125U
V_OS        85 31 2.99M
C30         21 22 15.92U  
R85         22 MID 30K NOISELESS  
R84         22 21 10K NOISELESS  
R83         21 MID 1 NOISELESS  
GVCCS10     24 MID 23 MID  -1
C29         25 MID 19.89F  
R82         23 25 10K NOISELESS  
R81         23 26 70k NOISELESS   
R80         26 MID 1 NOISELESS  
GVCCS9      26 MID 22 MID  -3.8
GVCCS4      21 MID CL_CLAMP 27  -87
R79         28 MID 1 NOISELESS  
XU1         29 MID MID 28 VCCS_LIM_ZO_0
R78         29 MID 101  NOISELESS  
C22         29 24 15.92F 
R65         29 24 10K NOISELESS  
R64         24 MID 1 NOISELESS  
R63         27 28 400k  NOISELESS  
XCLAWn      MID VIMON VEE_B 30 VCCS_LIM_CLAW-_0
Xe_n        ESDp 31 VNSE_0
Xi_nn       ESDn MID FEMT_0_0
Xi_np       MID 31 FEMT_0_0
S5          VEE ESDp VEE ESDp  S_VSWITCH_1
S4          VEE ESDn VEE ESDn  S_VSWITCH_2
S2          ESDn VCC ESDn VCC  S_VSWITCH_3
S3          ESDp VCC ESDp VCC  S_VSWITCH_4
C28         32 MID 1P 
R77         33 32 100  NOISELESS  
C27         34 MID 1P 
R76         35 34 100  NOISELESS  
R75         MID 36 1 NOISELESS  
GVCCS8      36 MID 37 MID  -1
R74         38 MID 1 NOISELESS  
GVCCS7      38 MID 39 MID  -1
C25         40 MID 25F 
R69         MID 40 1MEG  NOISELESS  
GVCCS6      40 MID VSENSE MID  -1U
C20         CLAMP MID 151.6N 
R68         MID CLAMP 1MEG  NOISELESS  
XVCCS_LIM_2 41 MID MID CLAMP VCCS_LIM_2_0
R44         MID 41 1MEG  NOISELESS  
XVCCS_LIM_1 42 43 MID 41 VCCS_LIM_1_0
Rdummy      MID 27 40k  NOISELESS  
R61         MID 44 273.3609  NOISELESS   
C16         44 45 1.1018N 
R58         45 44 100MEG   NOISELESS  
GVCCS2      45 MID VEE_B MID  -258.98M
R57         MID 45 1 NOISELESS  
R56         MID 46 273.3609  NOISELESS   
C15         46 47 1.1018N 
R55         47 46 100MEG   NOISELESS  
GVCCS1      47 MID VCC_B MID  -258.98M
R54         MID 47 1 NOISELESS  
R49         MID 48 337.4K   NOISELESS   
C14         48 49 591.7F 
R48         49 48 100MEG   NOISELESS  
G_adjust    49 MID ESDp MID  -44.81M
Rsrc        MID 49 1 NOISELESS  
XIQPos      VIMON MID MID VCC VCCS_LIMIT_IQ_0
XIQNeg      MID VIMON VEE MID VCCS_LIMIT_IQ_0
C_DIFF      ESDp ESDn 2P 
XCL_AMP     50 51 VIMON MID 52 53 CLAMP_AMP_LO_0
SOR_SWp     CLAMP 54 CLAMP 54  S_VSWITCH_5
SOR_SWn     55 CLAMP 55 CLAMP  S_VSWITCH_6
XGR_AMP     56 57 58 MID 59 60 CLAMP_AMP_HI_0
R39         56 MID 1t   NOISELESS   
R37         57 MID 1t   NOISELESS   
R42         VSENSE 58 1m   NOISELESS  
C19         58 MID 1F 
R38         59 MID 1 NOISELESS  
R36         MID 60 1 NOISELESS  
R40         59 61 1m   NOISELESS  
R41         60 62 1m   NOISELESS  
C17         61 MID 1F 
C18         MID 62 1F 
XGR_SRC     61 62 CLAMP MID VCCS_LIM_GR_0
R21         52 MID 1 NOISELESS  
R20         MID 53 1 NOISELESS  
R29         52 63 1m   NOISELESS  
R30         53 64 1m   NOISELESS  
C9          63 MID 1F 
C8          MID 64 1F 
XCL_SRC     63 64 CL_CLAMP MID VCCS_LIM_4_0
R22         50 MID 1t   NOISELESS   
R19         MID 51 1t   NOISELESS   
XCLAWp      VIMON MID 65 VCC_B VCCS_LIM_CLAW+_0
R12         65 VCC_B 1k   NOISELESS  
R16         65 66 1m   NOISELESS  
R13         VEE_B 30 1k   NOISELESS  
R17         67 30 1m   NOISELESS  
C6          67 MID 1F 
C5          MID 66 1F 
G2          VCC_CLP MID 66 MID  -1M
R15         VCC_CLP MID 1k   NOISELESS  
G3          VEE_CLP MID 67 MID  -1M
R14         MID VEE_CLP 1k   NOISELESS  
XCLAW_AMP   VCC_CLP VEE_CLP VOUT_S MID 68 69 CLAMP_AMP_LO_0
R26         VCC_CLP MID 1t   NOISELESS   
R23         VEE_CLP MID 1t   NOISELESS   
R25         68 MID 1 NOISELESS  
R24         MID 69 1 NOISELESS  
R27         68 70 1m   NOISELESS  
R28         69 71 1m   NOISELESS  
C11         70 MID 1F 
C10         MID 71 1F 
XCLAW_SRC   70 71 CLAW_CLAMP MID VCCS_LIM_3_0
H2          35 MID V11 -1
H3          33 MID V12 1
C12         SW_OL MID 100P 
R32         72 SW_OL 100  NOISELESS  
R31         72 MID 1 NOISELESS  
XOL_SENSE   MID 72 34 32 OL_SENSE_0
S1          21 22 SW_OL MID  S_VSWITCH_7
H1          73 MID V4 1K
S7          VEE OUT VEE OUT  S_VSWITCH_8
S6          OUT VCC OUT VCC  S_VSWITCH_9
R11         MID 74 1t   NOISELESS   
R18         74 VOUT_S 100  NOISELESS  
C7          VOUT_S MID 1P 
E5          74 MID OUT MID  1
C13         VIMON MID 1N 
R33         73 VIMON 100  NOISELESS  
R10         MID 73 1t   NOISELESS   
R47         75 VCLP 100  NOISELESS  
C24         VCLP MID 100P 
E4          75 MID CL_CLAMP MID  1
R46         MID CL_CLAMP 1k   NOISELESS  
G9          CL_CLAMP MID CLAW_CLAMP MID  -1M
R45         MID CLAW_CLAMP 1k   NOISELESS  
G8          CLAW_CLAMP MID 40 MID  -1M
R43         MID VSENSE 1k   NOISELESS  
G15         VSENSE MID CLAMP MID  -1M
C4          42 MID 1F 
R9          42 76 1m   NOISELESS  
R7          MID 77 1t   NOISELESS   
R6          78 MID 1t   NOISELESS   
R8          MID 76 1 NOISELESS  
XVCM_CLAMP  79 MID 76 MID 78 77 VCCS_EXT_LIM_0
E1          MID 0 80 0  1
R89         VEE_B 0 1 NOISELESS  
R5          81 VEE_B 1m   NOISELESS  
C3          81 0 1F 
R60         80 81 1MEG  NOISELESS  
C1          80 0 1 
R3          80 0 1t   NOISELESS   
R59         82 80 1MEG  NOISELESS  
C2          82 0 1F 
R4          VCC_B 82 1m   NOISELESS  
R88         VCC_B 0 1 NOISELESS  
G17         VEE_B 0 VEE 0  -1
G16         VCC_B 0 VCC 0  -1
R_PSR       83 79 1k   NOISELESS  
G_PSR       79 83 46 44  -1M
R2          43 ESDn 1m   NOISELESS  
R1          83 84 1m   NOISELESS  
R_CMR       85 84 1k   NOISELESS  
G_CMR       84 85 48 MID  -1M
C_CMn       ESDn MID 5.5P 
C_CMp       MID ESDp 5.5P 
R53         ESDn MID 1t   NOISELESS   
R52         MID ESDp 1t   NOISELESS   
R35         IN- ESDn 10m   NOISELESS  
R34         IN+ ESDp 10m   NOISELESS  

.MODEL S_VSWITCH_1 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_2 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_3 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_4 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_5 VSWITCH (RON=10M ROFF=1T VON=10M VOFF=0)
.MODEL S_VSWITCH_6 VSWITCH (RON=10M ROFF=1T VON=10M VOFF=0)
.MODEL S_VSWITCH_7 VSWITCH (RON=1M ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_8 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_9 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)

.ENDS LM324LV
*
.SUBCKT VCCS_LIM_ZO_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 100
.PARAM IPOS = 32E3
.PARAM INEG = -32E3
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*

.SUBCKT VCCS_LIM_CLAW-_0  VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {ABS(V(VC+,VC-))} =
+(00.0000, 0.00001)
+(14.0000, 0.000379)
+(28.0000, 0.000877)
+(37.3333, 0.001382)
+(37.8000, 0.00142)
+(38.7333, 0.001493)
+(39.6667, 0.001583)
+(40.6000, 0.001703)
+(41.5333, 0.00191)
+(42.0000, 0.00204)
.ENDS VCCS_LIM_CLAW-_0 
*

.SUBCKT VNSE_0  1 2
.PARAM FLW=10
.PARAM NLF=115
.PARAM NVR=27
.PARAM GLF={PWR(FLW,0.25)*NLF/1164}
.PARAM RNV={1.184*PWR(NVR,2)}
.MODEL DVN D KF={PWR(FLW,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVN
D2 8 0 DVN
E1 3 6 7 8 {GLF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNV}
R5 5 0 {RNV}
R6 3 4 1E9
R7 4 0 1E9
E3 1 2 3 4 1
.ENDS
*

.SUBCKT FEMT_0_0   1 2
.PARAM FLWF=0.001
.PARAM NLFF=23
.PARAM NVRF=23
.PARAM GLFF={PWR(FLWF,0.25)*NLFF/1164}
.PARAM RNVF={1.184*PWR(NVRF,2)}
.MODEL DVNF D KF={PWR(FLWF,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVNF
D2 8 0 DVNF
E1 3 6 7 8 {GLFF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNVF}
R5 5 0 {RNVF}
R6 3 4 1E9
R7 4 0 1E9
G1 1 2 3 4 1E-6
.ENDS
*

.SUBCKT VCCS_LIM_2_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 11.15E-3
.PARAM IPOS = 0.263
.PARAM INEG = -0.263
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*

.SUBCKT VCCS_LIM_1_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1E-4
.PARAM IPOS = .5
.PARAM INEG = -.5
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*

.SUBCKT VCCS_LIMIT_IQ_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1E-3
G1 IOUT- IOUT+ VALUE={IF( (V(VC+,VC-)<=0),0,GAIN*V(VC+,VC-) )}
.ENDS
*

.SUBCKT CLAMP_AMP_LO_0  VC+ VC- VIN COM VO+ VO-
.PARAM G=1
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS
*

.SUBCKT CLAMP_AMP_HI_0  VC+ VC- VIN COM VO+ VO-
.PARAM G=10
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS
*

.SUBCKT VCCS_LIM_GR_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 0.55
.PARAM INEG = -0.55
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*

.SUBCKT VCCS_LIM_4_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 1.122
.PARAM INEG = -1.122
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*

.SUBCKT VCCS_LIM_CLAW+_0  VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {ABS(V(VC+,VC-))} =
+(00.00, 0.000010)
+(13.67, 0.0003467)
+(27.33, 0.0007994)
+(36.44, 0.001309)
+(36.90, 0.001351)
+(37.81, 0.001455)
+(38.72, 0.001600)
+(39.63, 0.001812)
+(40.54, 0.002117)
+(41.00, 0.002292)
.ENDS VCCS_LIM_CLAW+_0 
*

.SUBCKT VCCS_LIM_3_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 0.47
.PARAM INEG = -0.47
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*

.SUBCKT OL_SENSE_0  COM SW+ OLN  OLP
GSW+ COM SW+ VALUE = {IF((V(OLN,COM)>10E-3 | V(OLP,COM)>10E-3),1,0)}
.ENDS
*

.SUBCKT VCCS_EXT_LIM_0  VIN+ VIN- IOUT- IOUT+ VP+ VP-
.PARAM GAIN = 1
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VIN+,VIN-),V(VP-,VIN-), V(VP+,VIN-))}
.ENDS
*

.subckt LM321LV IN+ IN- VCC VEE OUT
X IN+ IN- VCC VEE OUT LM324LV
.ends

.subckt LM358LV IN+ IN- VCC VEE OUT
X IN+ IN- VCC VEE OUT LM324LV
.ends