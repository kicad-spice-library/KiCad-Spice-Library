.MODEL 32ctq030h d
+IS=1e-15 RS=0.01 N=0.5 EG=1.07785
+XTI=4 BV=30 IBV=0.00175 CJO=2.11811e-09
+VJ=1.5 M=0.499425 FC=0.5 TT=0
+KF=0 AF=1
* Model generated on May 28, 96
* Model format: SPICE3

