* Version 2.0 Copyright � Linear Technology Corp. 10/19/04. All rights reserved.
*
* NODES 1 AND 8 = COMPENSATION PINS
*
.SUBCKT LM308 3 2 7 4 6 1 8
* USE C=30 PF IN MAIN CIRCUIT (CA TO CB).
* INPUT
RC1 7 80 8.842E+03
RC2 7 90 8.842E+03
Q1 80 2 10 QM1
Q2 90 3 11 QM2
DDM1 2 3 DM2
DDM2 3 2 DM2
C1 80 90 5.460E-12
RE1 10 12 2.245E+02
RE2 11 12 2.245E+02
IEE 12 4 6.003E-06
RE 12 0 3.332E+07
CE 12 0 1.579E-12
* INTERMEDIATE
GCM 0 8 12 0 1.131E-09
GA 8 0 80 90 1.131E-04
R2 8 0 1.000E+05
* EXTERNAL COMP CAP USED FOR C2 (SEE NOTE ABOVE).
GB 1 0 8 0 3.146E+01
* OUTPUT
RO1 1 6 1.111E+02
RO2 1 0 8.889E+02
RC 17 0 3.533E-04
GC 0 17 6 0 2.830E+03
D1 1 17 DM1
D2 17 1 DM1
D3 6 13 DM2
D4 14 6 DM2
VC 7 13 1.766E+00
VE 14 4 1.766E+00
IP 7 4 2.940E-04
DSUB 4 7 DM2
* MODELS
.MODEL QM1 NPN (IS=8.000E-16 BF=1.875E+03)
.MODEL QM2 NPN (IS=8.643E-16 BF=2.143E+03)
.MODEL DM1 D (IS=1.192E-10)
.MODEL DM2 D (IS=8.000E-16)
.ENDS LM308

