* AD633 LT Spice - a simplified MODEL of
* CONNECTIONS:
*                 Y2 -_   _- Vee
*               Y1 -_  | |  _- Z
*             X2 -_  | | | |  _- W
*           X1 -_  | | | | | | _- Vcc
*                | | | | | | | |
.SUBCKT AD633AN  1 2 3 4 5 6 7 8
*
R0   99    0    1Meg
R1   99    5    2Meg
R2   99    8    2Meg
R3   33   66    2k7
R4   66   99    300
B3   33   99    V={V(1,2)*V(3,4)}
R5   88   99    3k
B5   88   99    V={V(6,5)+I(R4)*300}
B4	  7	   5	V={if(V(88,99)>V(8,5),V(8,5),if(V(88,99)<0,0,V(88,99)))}
R95	 99    1    .1G
R96  99    2    .1G
R97  99    3    .1G
R98  99    4    .1G
R99  99    6    .1G
.ENDS
