test circuit #1 for pz analysis:high pass filter
r1 1 0 1k
r2 2 0 1k
c1 1 2 1.0e-12
.pz 1 0 2 0 cur pz
.print pz all
.end
