* 74HCT595.CIR
.subckt 74HCT595 DS SHCP _MR STCP _OE Q0 Q1 Q2 Q3 Q4 Q5 Q6 Q7 Q7S
.param Vdd=5
A1  DS  0 0 0 0 0 1 0 SCHMITT Vhigh={Vdd} tripdt=5n Vt=1.4 Vh=0.1
A2 SHCP 0 0 0 0 0 2 0 SCHMITT Vhigh={Vdd} tripdt=5n Vt=1.4 Vh=0.1
A3 _MR  0 0 0 0 3 0 0 SCHMITT Vhigh={Vdd} tripdt=5n Vt=1.4 Vh=0.1
A4 STCP 0 0 0 0 0 4 0 SCHMITT Vhigh={Vdd} tripdt=5n Vt=1.4 Vh=0.1
A5 _OE 0 0 0 0 OE 0 0 SCHMITT Vhigh={Vdd} tripdt=5n Vt=1.4 Vh=0.1
A6   1 0 2 0 3 0  5 0 DFLOP Vhigh={Vdd} td=10n tripdt=5n
A7   5 0 2 0 3 0  6 0 DFLOP Vhigh={Vdd} td=10n tripdt=5n
A8   6 0 2 0 3 0  7 0 DFLOP Vhigh={Vdd} td=10n tripdt=5n
A9   7 0 2 0 3 0  8 0 DFLOP Vhigh={Vdd} td=10n tripdt=5n
A10  8 0 2 0 3 0  9 0 DFLOP Vhigh={Vdd} td=10n tripdt=5n
A11  9 0 2 0 3 0 10 0 DFLOP Vhigh={Vdd} td=10n tripdt=5n
A12 10 0 2 0 3 0 11 0 DFLOP Vhigh={Vdd} td=10n tripdt=5n
A13 11 0 2 0 3 0 Q7S 0 DFLOP Vhigh={Vdd} td=10n tripdt=5n Rout=50
A14  5 0 4 0 0 0 12 0 DFLOP Vhigh={Vdd} td=10n tripdt=5n
A15  6 0 4 0 0 0 13 0 DFLOP Vhigh={Vdd} td=10n tripdt=5n
A16  7 0 4 0 0 0 14 0 DFLOP Vhigh={Vdd} td=10n tripdt=5n
A17  8 0 4 0 0 0 15 0 DFLOP Vhigh={Vdd} td=10n tripdt=5n
A18  9 0 4 0 0 0 16 0 DFLOP Vhigh={Vdd} td=10n tripdt=5n
A19 10 0 4 0 0 0 17 0 DFLOP Vhigh={Vdd} td=10n tripdt=5n
A20 11 0 4 0 0 0 18 0 DFLOP Vhigh={Vdd} td=10n tripdt=5n
A21 Q7S 0 4 0 0 0 19 0 DFLOP Vhigh={Vdd} td=10n tripdt=5n
.func tri(x)=inv(x)*1G+30
R1  6 Q0 R=tri(V(OE))
R2  8 Q1 R=tri(V(OE))
R3 10 Q2 R=tri(V(OE))
R4 12 Q3 R=tri(V(OE))
R5 14 Q4 R=tri(V(OE))
R6 16 Q5 R=tri(V(OE))
R7 18 Q6 R=tri(V(OE))
R8 19 Q7 R=tri(V(OE))
.ends 74HCT595
