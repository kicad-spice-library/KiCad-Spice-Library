.MODEL 10bq015 d
+IS=1.66692e-05 RS=0.0549971 N=1.0339 EG=0.6
+XTI=0.5 BV=15 IBV=0.001 CJO=4.70891e-10
+VJ=1.5 M=0.699718 FC=0.5 TT=0
+KF=0 AF=1
* Model generated on May 28, 96
* Model format: SPICE3

