.MODEL 20clq045 d
+IS=5.55194e-10 RS=0.01 N=0.736126 EG=0.6
+XTI=0.5 BV=45 IBV=0.005 CJO=2.42073e-09
+VJ=0.470122 M=0.477502 FC=0.5 TT=0
+KF=0 AF=1
* Model generated on May 28, 96
* Model format: SPICE3

