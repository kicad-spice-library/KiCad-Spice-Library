.MODEL 20ets12avg d
+IS=3.14987e-10 RS=0.01 N=1.37516 EG=1.06967
+XTI=4 BV=1200 IBV=0.0001 CJO=1e-11
+VJ=0.7 M=0.5 FC=0.5 TT=1e-09
+KF=0 AF=1
* Model generated on Apr 26, 96
* Model format: SPICE3

