BJT Characteristics

*.lib bipolar.lib

.MODEL BC107BP NPN IS=1.8E-14 ISE=5.0E-14 NF=.9955 NE=1.46 BF=220 BR=35.5
+IKF=.14 IKR=.03 ISC=1.72E-13 NC=1.27 NR=1.005 RB=.56 RE=.6 RC=0.25 VAF=80
+VAR=12.5 CJE=13E-12 TF=.64E-9 CJC=4E-12 TR=50.72E-9 VJC=.54 MJC=.33

.model BC107    NPN(Is=1.527f Xti=3 Eg=1.11 Vaf=106.8 Bf=334.5 Ne=1.642
+               Ise=222f Ikf=.1596 Xtb=1.5 Br=.788 Nc=2 Isc=0 Ikr=0 Re=.6 Rc=0.25
+               Cjc=6.072p Mjc=.3333 Vjc=.75 Fc=.5 Cje=10.67p Mje=.3333 Vje=.75
+               Tr=10n Tf=471.8p Itf=0 Vtf=0 Xtf=0)

* Circuit to plot curves of Ic versus Vce for comparison with a datasheet

Ib 0 1 DC 50e-6
Q1 2 1 0 BC107
Vce 2 0 0V

.control
destroy all
save all
foreach basecurrent 50e-6 100e-6 200e-6 300e-6 500e-6 750e-6 1000e-6
    alter @Ib[DC] = $basecurrent
    dc Vce 0 4 0.1
end

plot abs(dc1.vce#branch)
+ abs(dc2.vce#branch)
+ abs(dc3.vce#branch)
+ abs(dc4.vce#branch)
+ abs(dc5.vce#branch)
+ xlabel Vce
+ ylabel Ic

.endc
